Schema_Prototype

.option savecurrents
.option interp
.OP
*.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END